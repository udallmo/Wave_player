// QD1.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module QD1 (
		inout  wire        audio_i2c_SDAT,              //      audio_i2c.SDAT
		output wire        audio_i2c_SCLK,              //               .SCLK
		output wire        audio_mclk_clk,              //     audio_mclk.clk
		input  wire        audio_out_ADCDAT,            //      audio_out.ADCDAT
		input  wire        audio_out_ADCLRCK,           //               .ADCLRCK
		input  wire        audio_out_BCLK,              //               .BCLK
		output wire        audio_out_DACDAT,            //               .DACDAT
		input  wire        audio_out_DACLRCK,           //               .DACLRCK
		input  wire [3:0]  button_pio_export,           //     button_pio.export
		input  wire        clk_50_clk,                  //         clk_50.clk
		output wire [7:0]  dual_7_segment_segment_data, // dual_7_segment.segment_data
		output wire        dual_7_segment_digit1,       //               .digit1
		output wire        dual_7_segment_digit2,       //               .digit2
		output wire        egm_interface_stimulus,      //  egm_interface.stimulus
		input  wire        egm_interface_response,      //               .response
		output wire [3:0]  egm_interface_egm_leds,      //               .egm_leds
		output wire        lcd_display_RS,              //    lcd_display.RS
		output wire        lcd_display_RW,              //               .RW
		inout  wire [7:0]  lcd_display_data,            //               .data
		output wire        lcd_display_E,               //               .E
		output wire [3:0]  led_pio_export,              //        led_pio.export
		input  wire        reset_reset_n,               //          reset.reset_n
		output wire        response_out_export,         //   response_out.export
		output wire [11:0] sdram_0_addr,                //        sdram_0.addr
		output wire [1:0]  sdram_0_ba,                  //               .ba
		output wire        sdram_0_cas_n,               //               .cas_n
		output wire        sdram_0_cke,                 //               .cke
		output wire        sdram_0_cs_n,                //               .cs_n
		inout  wire [15:0] sdram_0_dq,                  //               .dq
		output wire [1:0]  sdram_0_dqm,                 //               .dqm
		output wire        sdram_0_ras_n,               //               .ras_n
		output wire        sdram_0_we_n,                //               .we_n
		output wire        sdram_clk_clk,               //      sdram_clk.clk
		output wire        spi_master_cs,               //     spi_master.cs
		output wire        spi_master_sclk,             //               .sclk
		output wire        spi_master_mosi,             //               .mosi
		input  wire        spi_master_miso,             //               .miso
		input  wire        spi_master_cd,               //               .cd
		input  wire        spi_master_wp,               //               .wp
		input  wire        stimulus_in_export,          //    stimulus_in.export
		input  wire [7:0]  switch_pio_export,           //     switch_pio.export
		input  wire        uart_rxd,                    //           uart.rxd
		output wire        uart_txd                     //               .txd
	);

	wire         altpll_0_c2_clk;                                                       // altpll_0:c2 -> [Audio:clk, audio_i2c_config:clk, button_pio:clk, egm:clk, irq_mapper:clk, jtag_uart_0:clk, lcd_display:clk, led_pio:clk, mm_interconnect_0:altpll_0_c2_clk, nios2_gen2_0:clk, response_out:clk, rst_controller:clk, sdram_0:clk, seven_seg_pio:clk, spi_master:clk, stimulus_in:clk, switch_pio:clk, sysid_qsys_0:clock, system_timer:clk, timer_0:clk, uart:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                     // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                  // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                  // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [24:0] nios2_gen2_0_data_master_address;                                      // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                   // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                         // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                                // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                                        // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                    // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                              // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                           // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [24:0] nios2_gen2_0_instruction_master_address;                               // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                  // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                         // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_audio_avalon_audio_slave_chipselect;                 // mm_interconnect_0:Audio_avalon_audio_slave_chipselect -> Audio:chipselect
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_readdata;                   // Audio:readdata -> mm_interconnect_0:Audio_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_avalon_audio_slave_address;                    // mm_interconnect_0:Audio_avalon_audio_slave_address -> Audio:address
	wire         mm_interconnect_0_audio_avalon_audio_slave_read;                       // mm_interconnect_0:Audio_avalon_audio_slave_read -> Audio:read
	wire         mm_interconnect_0_audio_avalon_audio_slave_write;                      // mm_interconnect_0:Audio_avalon_audio_slave_write -> Audio:write
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_writedata;                  // mm_interconnect_0:Audio_avalon_audio_slave_writedata -> Audio:writedata
	wire  [31:0] mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_readdata;    // audio_i2c_config:readdata -> mm_interconnect_0:audio_i2c_config_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_waitrequest; // audio_i2c_config:waitrequest -> mm_interconnect_0:audio_i2c_config_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_address;     // mm_interconnect_0:audio_i2c_config_avalon_av_config_slave_address -> audio_i2c_config:address
	wire         mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_read;        // mm_interconnect_0:audio_i2c_config_avalon_av_config_slave_read -> audio_i2c_config:read
	wire   [3:0] mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_byteenable;  // mm_interconnect_0:audio_i2c_config_avalon_av_config_slave_byteenable -> audio_i2c_config:byteenable
	wire         mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_write;       // mm_interconnect_0:audio_i2c_config_avalon_av_config_slave_write -> audio_i2c_config:write
	wire  [31:0] mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_writedata;   // mm_interconnect_0:audio_i2c_config_avalon_av_config_slave_writedata -> audio_i2c_config:writedata
	wire         mm_interconnect_0_egm_avalon_egm_slave_chipselect;                     // mm_interconnect_0:egm_avalon_egm_slave_chipselect -> egm:chipselect
	wire  [31:0] mm_interconnect_0_egm_avalon_egm_slave_readdata;                       // egm:readdata -> mm_interconnect_0:egm_avalon_egm_slave_readdata
	wire   [2:0] mm_interconnect_0_egm_avalon_egm_slave_address;                        // mm_interconnect_0:egm_avalon_egm_slave_address -> egm:address
	wire         mm_interconnect_0_egm_avalon_egm_slave_read;                           // mm_interconnect_0:egm_avalon_egm_slave_read -> egm:read
	wire         mm_interconnect_0_egm_avalon_egm_slave_write;                          // mm_interconnect_0:egm_avalon_egm_slave_write -> egm:write
	wire  [31:0] mm_interconnect_0_egm_avalon_egm_slave_writedata;                      // mm_interconnect_0:egm_avalon_egm_slave_writedata -> egm:writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;            // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;              // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;           // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;               // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                 // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;             // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_seven_seg_pio_avalon_slave_0_chipselect;             // mm_interconnect_0:seven_seg_pio_avalon_slave_0_chipselect -> seven_seg_pio:chipselect
	wire  [31:0] mm_interconnect_0_seven_seg_pio_avalon_slave_0_readdata;               // seven_seg_pio:readdata -> mm_interconnect_0:seven_seg_pio_avalon_slave_0_readdata
	wire   [2:0] mm_interconnect_0_seven_seg_pio_avalon_slave_0_address;                // mm_interconnect_0:seven_seg_pio_avalon_slave_0_address -> seven_seg_pio:address
	wire         mm_interconnect_0_seven_seg_pio_avalon_slave_0_read;                   // mm_interconnect_0:seven_seg_pio_avalon_slave_0_read -> seven_seg_pio:read
	wire         mm_interconnect_0_seven_seg_pio_avalon_slave_0_write;                  // mm_interconnect_0:seven_seg_pio_avalon_slave_0_write -> seven_seg_pio:write
	wire  [31:0] mm_interconnect_0_seven_seg_pio_avalon_slave_0_writedata;              // mm_interconnect_0:seven_seg_pio_avalon_slave_0_writedata -> seven_seg_pio:writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                 // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                  // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire   [7:0] mm_interconnect_0_lcd_display_control_slave_readdata;                  // lcd_display:readdata -> mm_interconnect_0:lcd_display_control_slave_readdata
	wire   [1:0] mm_interconnect_0_lcd_display_control_slave_address;                   // mm_interconnect_0:lcd_display_control_slave_address -> lcd_display:address
	wire         mm_interconnect_0_lcd_display_control_slave_read;                      // mm_interconnect_0:lcd_display_control_slave_read -> lcd_display:read
	wire         mm_interconnect_0_lcd_display_control_slave_begintransfer;             // mm_interconnect_0:lcd_display_control_slave_begintransfer -> lcd_display:begintransfer
	wire         mm_interconnect_0_lcd_display_control_slave_write;                     // mm_interconnect_0:lcd_display_control_slave_write -> lcd_display:write
	wire   [7:0] mm_interconnect_0_lcd_display_control_slave_writedata;                 // mm_interconnect_0:lcd_display_control_slave_writedata -> lcd_display:writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;               // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;            // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;             // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_0_s1_chipselect;                               // mm_interconnect_0:sdram_0_s1_chipselect -> sdram_0:az_cs
	wire  [15:0] mm_interconnect_0_sdram_0_s1_readdata;                                 // sdram_0:za_data -> mm_interconnect_0:sdram_0_s1_readdata
	wire         mm_interconnect_0_sdram_0_s1_waitrequest;                              // sdram_0:za_waitrequest -> mm_interconnect_0:sdram_0_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_0_s1_address;                                  // mm_interconnect_0:sdram_0_s1_address -> sdram_0:az_addr
	wire         mm_interconnect_0_sdram_0_s1_read;                                     // mm_interconnect_0:sdram_0_s1_read -> sdram_0:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_0_s1_byteenable;                               // mm_interconnect_0:sdram_0_s1_byteenable -> sdram_0:az_be_n
	wire         mm_interconnect_0_sdram_0_s1_readdatavalid;                            // sdram_0:za_valid -> mm_interconnect_0:sdram_0_s1_readdatavalid
	wire         mm_interconnect_0_sdram_0_s1_write;                                    // mm_interconnect_0:sdram_0_s1_write -> sdram_0:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_0_s1_writedata;                                // mm_interconnect_0:sdram_0_s1_writedata -> sdram_0:az_data
	wire         mm_interconnect_0_led_pio_s1_chipselect;                               // mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_0_led_pio_s1_readdata;                                 // led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_led_pio_s1_address;                                  // mm_interconnect_0:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_0_led_pio_s1_write;                                    // mm_interconnect_0:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_0_led_pio_s1_writedata;                                // mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	wire         mm_interconnect_0_button_pio_s1_chipselect;                            // mm_interconnect_0:button_pio_s1_chipselect -> button_pio:chipselect
	wire  [31:0] mm_interconnect_0_button_pio_s1_readdata;                              // button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_button_pio_s1_address;                               // mm_interconnect_0:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_0_button_pio_s1_write;                                 // mm_interconnect_0:button_pio_s1_write -> button_pio:write_n
	wire  [31:0] mm_interconnect_0_button_pio_s1_writedata;                             // mm_interconnect_0:button_pio_s1_writedata -> button_pio:writedata
	wire  [31:0] mm_interconnect_0_switch_pio_s1_readdata;                              // switch_pio:readdata -> mm_interconnect_0:switch_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_switch_pio_s1_address;                               // mm_interconnect_0:switch_pio_s1_address -> switch_pio:address
	wire         mm_interconnect_0_uart_s1_chipselect;                                  // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                                    // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                                     // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                                        // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                               // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                                       // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                                   // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_system_timer_s1_chipselect;                          // mm_interconnect_0:system_timer_s1_chipselect -> system_timer:chipselect
	wire  [15:0] mm_interconnect_0_system_timer_s1_readdata;                            // system_timer:readdata -> mm_interconnect_0:system_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_system_timer_s1_address;                             // mm_interconnect_0:system_timer_s1_address -> system_timer:address
	wire         mm_interconnect_0_system_timer_s1_write;                               // mm_interconnect_0:system_timer_s1_write -> system_timer:write_n
	wire  [15:0] mm_interconnect_0_system_timer_s1_writedata;                           // mm_interconnect_0:system_timer_s1_writedata -> system_timer:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                               // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                                 // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                  // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                    // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                                // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_spi_master_s1_chipselect;                            // mm_interconnect_0:spi_master_s1_chipselect -> spi_master:chipselect
	wire  [31:0] mm_interconnect_0_spi_master_s1_readdata;                              // spi_master:readdata -> mm_interconnect_0:spi_master_s1_readdata
	wire   [2:0] mm_interconnect_0_spi_master_s1_address;                               // mm_interconnect_0:spi_master_s1_address -> spi_master:address
	wire         mm_interconnect_0_spi_master_s1_read;                                  // mm_interconnect_0:spi_master_s1_read -> spi_master:read
	wire         mm_interconnect_0_spi_master_s1_write;                                 // mm_interconnect_0:spi_master_s1_write -> spi_master:write
	wire  [31:0] mm_interconnect_0_spi_master_s1_writedata;                             // mm_interconnect_0:spi_master_s1_writedata -> spi_master:writedata
	wire         mm_interconnect_0_response_out_s1_chipselect;                          // mm_interconnect_0:response_out_s1_chipselect -> response_out:chipselect
	wire  [31:0] mm_interconnect_0_response_out_s1_readdata;                            // response_out:readdata -> mm_interconnect_0:response_out_s1_readdata
	wire   [1:0] mm_interconnect_0_response_out_s1_address;                             // mm_interconnect_0:response_out_s1_address -> response_out:address
	wire         mm_interconnect_0_response_out_s1_write;                               // mm_interconnect_0:response_out_s1_write -> response_out:write_n
	wire  [31:0] mm_interconnect_0_response_out_s1_writedata;                           // mm_interconnect_0:response_out_s1_writedata -> response_out:writedata
	wire         mm_interconnect_0_stimulus_in_s1_chipselect;                           // mm_interconnect_0:stimulus_in_s1_chipselect -> stimulus_in:chipselect
	wire  [31:0] mm_interconnect_0_stimulus_in_s1_readdata;                             // stimulus_in:readdata -> mm_interconnect_0:stimulus_in_s1_readdata
	wire   [1:0] mm_interconnect_0_stimulus_in_s1_address;                              // mm_interconnect_0:stimulus_in_s1_address -> stimulus_in:address
	wire         mm_interconnect_0_stimulus_in_s1_write;                                // mm_interconnect_0:stimulus_in_s1_write -> stimulus_in:write_n
	wire  [31:0] mm_interconnect_0_stimulus_in_s1_writedata;                            // mm_interconnect_0:stimulus_in_s1_writedata -> stimulus_in:writedata
	wire         irq_mapper_receiver0_irq;                                              // Audio:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                              // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                              // uart:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                              // button_pio:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                              // system_timer:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                              // timer_0:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                              // stimulus_in:irq -> irq_mapper:receiver6_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                  // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                        // rst_controller:reset_out -> [Audio:reset, audio_i2c_config:reset, button_pio:reset_n, egm:reset, irq_mapper:reset, jtag_uart_0:rst_n, lcd_display:reset_n, led_pio:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, response_out:reset_n, rst_translator:in_reset, sdram_0:reset_n, seven_seg_pio:reset, spi_master:reset, stimulus_in:reset_n, switch_pio:reset_n, sysid_qsys_0:reset_n, system_timer:reset_n, timer_0:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                                    // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                    // rst_controller_001:reset_out -> altpll_0:reset

	QD1_Audio audio (
		.clk         (altpll_0_c2_clk),                                       //                clk.clk
		.reset       (rst_controller_reset_out_reset),                        //              reset.reset
		.address     (mm_interconnect_0_audio_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audio_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audio_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audio_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audio_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audio_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver0_irq),                              //          interrupt.irq
		.AUD_ADCDAT  (audio_out_ADCDAT),                                      // external_interface.export
		.AUD_ADCLRCK (audio_out_ADCLRCK),                                     //                   .export
		.AUD_BCLK    (audio_out_BCLK),                                        //                   .export
		.AUD_DACDAT  (audio_out_DACDAT),                                      //                   .export
		.AUD_DACLRCK (audio_out_DACLRCK)                                      //                   .export
	);

	QD1_altpll_0 altpll_0 (
		.clk       (clk_50_clk),                         //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (sdram_clk_clk),                      //                    c0.clk
		.c1        (audio_mclk_clk),                     //                    c1.clk
		.c2        (altpll_0_c2_clk),                    //                    c2.clk
		.areset    (),                                   //        areset_conduit.export
		.locked    (),                                   //        locked_conduit.export
		.phasedone ()                                    //     phasedone_conduit.export
	);

	QD1_audio_i2c_config audio_i2c_config (
		.clk         (altpll_0_c2_clk),                                                       //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                        //                  reset.reset
		.address     (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_i2c_SDAT),                                                        //     external_interface.export
		.I2C_SCLK    (audio_i2c_SCLK)                                                         //                       .export
	);

	QD1_button_pio button_pio (
		.clk        (altpll_0_c2_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                    //                 irq.irq
	);

	egm egm (
		.reset      (rst_controller_reset_out_reset),                    //            reset.reset
		.chipselect (mm_interconnect_0_egm_avalon_egm_slave_chipselect), // avalon_egm_slave.chipselect
		.address    (mm_interconnect_0_egm_avalon_egm_slave_address),    //                 .address
		.write      (mm_interconnect_0_egm_avalon_egm_slave_write),      //                 .write
		.writedata  (mm_interconnect_0_egm_avalon_egm_slave_writedata),  //                 .writedata
		.read       (mm_interconnect_0_egm_avalon_egm_slave_read),       //                 .read
		.readdata   (mm_interconnect_0_egm_avalon_egm_slave_readdata),   //                 .readdata
		.STIM       (egm_interface_stimulus),                            //        interface.stimulus
		.RESP       (egm_interface_response),                            //                 .response
		.EGM_LEDS   (egm_interface_egm_leds),                            //                 .egm_leds
		.clk        (altpll_0_c2_clk)                                    //              clk.clk
	);

	QD1_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c2_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	QD1_lcd_display lcd_display (
		.reset_n       (~rst_controller_reset_out_reset),                           //         reset.reset_n
		.clk           (altpll_0_c2_clk),                                           //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_display_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_display_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_display_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_display_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_display_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_display_control_slave_address),       //              .address
		.LCD_RS        (lcd_display_RS),                                            //      external.export
		.LCD_RW        (lcd_display_RW),                                            //              .export
		.LCD_data      (lcd_display_data),                                          //              .export
		.LCD_E         (lcd_display_E)                                              //              .export
	);

	QD1_led_pio led_pio (
		.clk        (altpll_0_c2_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_export)                           // external_connection.export
	);

	QD1_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (altpll_0_c2_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	QD1_response_out response_out (
		.clk        (altpll_0_c2_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_response_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_response_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_response_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_response_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_response_out_s1_readdata),   //                    .readdata
		.out_port   (response_out_export)                           // external_connection.export
	);

	QD1_sdram_0 sdram_0 (
		.clk            (altpll_0_c2_clk),                            //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),            // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_0_addr),                               //  wire.export
		.zs_ba          (sdram_0_ba),                                 //      .export
		.zs_cas_n       (sdram_0_cas_n),                              //      .export
		.zs_cke         (sdram_0_cke),                                //      .export
		.zs_cs_n        (sdram_0_cs_n),                               //      .export
		.zs_dq          (sdram_0_dq),                                 //      .export
		.zs_dqm         (sdram_0_dqm),                                //      .export
		.zs_ras_n       (sdram_0_ras_n),                              //      .export
		.zs_we_n        (sdram_0_we_n)                                //      .export
	);

	dual7segment seven_seg_pio (
		.chipselect (mm_interconnect_0_seven_seg_pio_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.address    (mm_interconnect_0_seven_seg_pio_avalon_slave_0_address),    //               .address
		.write      (mm_interconnect_0_seven_seg_pio_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_seven_seg_pio_avalon_slave_0_writedata),  //               .writedata
		.read       (mm_interconnect_0_seven_seg_pio_avalon_slave_0_read),       //               .read
		.readdata   (mm_interconnect_0_seven_seg_pio_avalon_slave_0_readdata),   //               .readdata
		.reset      (rst_controller_reset_out_reset),                            //          reset.reset
		.DOUT       (dual_7_segment_segment_data),                               // dual_7_segment.segment_data
		.DIG2       (dual_7_segment_digit1),                                     //               .digit1
		.DIG1       (dual_7_segment_digit2),                                     //               .digit2
		.clk        (altpll_0_c2_clk)                                            //            clk.clk
	);

	spi_master_if spi_master (
		.reset      (rst_controller_reset_out_reset),             //    reset.reset
		.clk        (altpll_0_c2_clk),                            //      clk.clk
		.chipselect (mm_interconnect_0_spi_master_s1_chipselect), //       s1.chipselect
		.address    (mm_interconnect_0_spi_master_s1_address),    //         .address
		.write      (mm_interconnect_0_spi_master_s1_write),      //         .write
		.writedata  (mm_interconnect_0_spi_master_s1_writedata),  //         .writedata
		.read       (mm_interconnect_0_spi_master_s1_read),       //         .read
		.readdata   (mm_interconnect_0_spi_master_s1_readdata),   //         .readdata
		.cs         (spi_master_cs),                              // external.export
		.sclk       (spi_master_sclk),                            //         .export
		.mosi       (spi_master_mosi),                            //         .export
		.miso       (spi_master_miso),                            //         .export
		.cd         (spi_master_cd),                              //         .export
		.wp         (spi_master_wp)                               //         .export
	);

	QD1_stimulus_in stimulus_in (
		.clk        (altpll_0_c2_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_stimulus_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_stimulus_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_stimulus_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_stimulus_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_stimulus_in_s1_readdata),   //                    .readdata
		.in_port    (stimulus_in_export),                          // external_connection.export
		.irq        (irq_mapper_receiver6_irq)                     //                 irq.irq
	);

	QD1_switch_pio switch_pio (
		.clk      (altpll_0_c2_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_switch_pio_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switch_pio_s1_readdata), //                    .readdata
		.in_port  (switch_pio_export)                         // external_connection.export
	);

	QD1_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c2_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	QD1_system_timer system_timer (
		.clk        (altpll_0_c2_clk),                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              // reset.reset_n
		.address    (mm_interconnect_0_system_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_system_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_system_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_system_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_system_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                      //   irq.irq
	);

	QD1_system_timer timer_0 (
		.clk        (altpll_0_c2_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                 //   irq.irq
	);

	QD1_uart uart (
		.clk           (altpll_0_c2_clk),                         //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.dataavailable (),                                        //                    .dataavailable
		.readyfordata  (),                                        //                    .readyfordata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	QD1_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c2_clk                                     (altpll_0_c2_clk),                                                       //                              altpll_0_c2.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                                        // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                    (nios2_gen2_0_data_master_address),                                      //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                (nios2_gen2_0_data_master_waitrequest),                                  //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable                 (nios2_gen2_0_data_master_byteenable),                                   //                                         .byteenable
		.nios2_gen2_0_data_master_read                       (nios2_gen2_0_data_master_read),                                         //                                         .read
		.nios2_gen2_0_data_master_readdata                   (nios2_gen2_0_data_master_readdata),                                     //                                         .readdata
		.nios2_gen2_0_data_master_readdatavalid              (nios2_gen2_0_data_master_readdatavalid),                                //                                         .readdatavalid
		.nios2_gen2_0_data_master_write                      (nios2_gen2_0_data_master_write),                                        //                                         .write
		.nios2_gen2_0_data_master_writedata                  (nios2_gen2_0_data_master_writedata),                                    //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess                (nios2_gen2_0_data_master_debugaccess),                                  //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address             (nios2_gen2_0_instruction_master_address),                               //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest         (nios2_gen2_0_instruction_master_waitrequest),                           //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read                (nios2_gen2_0_instruction_master_read),                                  //                                         .read
		.nios2_gen2_0_instruction_master_readdata            (nios2_gen2_0_instruction_master_readdata),                              //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid       (nios2_gen2_0_instruction_master_readdatavalid),                         //                                         .readdatavalid
		.Audio_avalon_audio_slave_address                    (mm_interconnect_0_audio_avalon_audio_slave_address),                    //                 Audio_avalon_audio_slave.address
		.Audio_avalon_audio_slave_write                      (mm_interconnect_0_audio_avalon_audio_slave_write),                      //                                         .write
		.Audio_avalon_audio_slave_read                       (mm_interconnect_0_audio_avalon_audio_slave_read),                       //                                         .read
		.Audio_avalon_audio_slave_readdata                   (mm_interconnect_0_audio_avalon_audio_slave_readdata),                   //                                         .readdata
		.Audio_avalon_audio_slave_writedata                  (mm_interconnect_0_audio_avalon_audio_slave_writedata),                  //                                         .writedata
		.Audio_avalon_audio_slave_chipselect                 (mm_interconnect_0_audio_avalon_audio_slave_chipselect),                 //                                         .chipselect
		.audio_i2c_config_avalon_av_config_slave_address     (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_address),     //  audio_i2c_config_avalon_av_config_slave.address
		.audio_i2c_config_avalon_av_config_slave_write       (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_write),       //                                         .write
		.audio_i2c_config_avalon_av_config_slave_read        (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_read),        //                                         .read
		.audio_i2c_config_avalon_av_config_slave_readdata    (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_readdata),    //                                         .readdata
		.audio_i2c_config_avalon_av_config_slave_writedata   (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_writedata),   //                                         .writedata
		.audio_i2c_config_avalon_av_config_slave_byteenable  (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_byteenable),  //                                         .byteenable
		.audio_i2c_config_avalon_av_config_slave_waitrequest (mm_interconnect_0_audio_i2c_config_avalon_av_config_slave_waitrequest), //                                         .waitrequest
		.button_pio_s1_address                               (mm_interconnect_0_button_pio_s1_address),                               //                            button_pio_s1.address
		.button_pio_s1_write                                 (mm_interconnect_0_button_pio_s1_write),                                 //                                         .write
		.button_pio_s1_readdata                              (mm_interconnect_0_button_pio_s1_readdata),                              //                                         .readdata
		.button_pio_s1_writedata                             (mm_interconnect_0_button_pio_s1_writedata),                             //                                         .writedata
		.button_pio_s1_chipselect                            (mm_interconnect_0_button_pio_s1_chipselect),                            //                                         .chipselect
		.egm_avalon_egm_slave_address                        (mm_interconnect_0_egm_avalon_egm_slave_address),                        //                     egm_avalon_egm_slave.address
		.egm_avalon_egm_slave_write                          (mm_interconnect_0_egm_avalon_egm_slave_write),                          //                                         .write
		.egm_avalon_egm_slave_read                           (mm_interconnect_0_egm_avalon_egm_slave_read),                           //                                         .read
		.egm_avalon_egm_slave_readdata                       (mm_interconnect_0_egm_avalon_egm_slave_readdata),                       //                                         .readdata
		.egm_avalon_egm_slave_writedata                      (mm_interconnect_0_egm_avalon_egm_slave_writedata),                      //                                         .writedata
		.egm_avalon_egm_slave_chipselect                     (mm_interconnect_0_egm_avalon_egm_slave_chipselect),                     //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),               //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                 //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                  //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),              //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),             //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),           //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),            //                                         .chipselect
		.lcd_display_control_slave_address                   (mm_interconnect_0_lcd_display_control_slave_address),                   //                lcd_display_control_slave.address
		.lcd_display_control_slave_write                     (mm_interconnect_0_lcd_display_control_slave_write),                     //                                         .write
		.lcd_display_control_slave_read                      (mm_interconnect_0_lcd_display_control_slave_read),                      //                                         .read
		.lcd_display_control_slave_readdata                  (mm_interconnect_0_lcd_display_control_slave_readdata),                  //                                         .readdata
		.lcd_display_control_slave_writedata                 (mm_interconnect_0_lcd_display_control_slave_writedata),                 //                                         .writedata
		.lcd_display_control_slave_begintransfer             (mm_interconnect_0_lcd_display_control_slave_begintransfer),             //                                         .begintransfer
		.led_pio_s1_address                                  (mm_interconnect_0_led_pio_s1_address),                                  //                               led_pio_s1.address
		.led_pio_s1_write                                    (mm_interconnect_0_led_pio_s1_write),                                    //                                         .write
		.led_pio_s1_readdata                                 (mm_interconnect_0_led_pio_s1_readdata),                                 //                                         .readdata
		.led_pio_s1_writedata                                (mm_interconnect_0_led_pio_s1_writedata),                                //                                         .writedata
		.led_pio_s1_chipselect                               (mm_interconnect_0_led_pio_s1_chipselect),                               //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),                //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                  //                                         .write
		.nios2_gen2_0_debug_mem_slave_read                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                   //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),               //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),              //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),             //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),            //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),            //                                         .debugaccess
		.response_out_s1_address                             (mm_interconnect_0_response_out_s1_address),                             //                          response_out_s1.address
		.response_out_s1_write                               (mm_interconnect_0_response_out_s1_write),                               //                                         .write
		.response_out_s1_readdata                            (mm_interconnect_0_response_out_s1_readdata),                            //                                         .readdata
		.response_out_s1_writedata                           (mm_interconnect_0_response_out_s1_writedata),                           //                                         .writedata
		.response_out_s1_chipselect                          (mm_interconnect_0_response_out_s1_chipselect),                          //                                         .chipselect
		.sdram_0_s1_address                                  (mm_interconnect_0_sdram_0_s1_address),                                  //                               sdram_0_s1.address
		.sdram_0_s1_write                                    (mm_interconnect_0_sdram_0_s1_write),                                    //                                         .write
		.sdram_0_s1_read                                     (mm_interconnect_0_sdram_0_s1_read),                                     //                                         .read
		.sdram_0_s1_readdata                                 (mm_interconnect_0_sdram_0_s1_readdata),                                 //                                         .readdata
		.sdram_0_s1_writedata                                (mm_interconnect_0_sdram_0_s1_writedata),                                //                                         .writedata
		.sdram_0_s1_byteenable                               (mm_interconnect_0_sdram_0_s1_byteenable),                               //                                         .byteenable
		.sdram_0_s1_readdatavalid                            (mm_interconnect_0_sdram_0_s1_readdatavalid),                            //                                         .readdatavalid
		.sdram_0_s1_waitrequest                              (mm_interconnect_0_sdram_0_s1_waitrequest),                              //                                         .waitrequest
		.sdram_0_s1_chipselect                               (mm_interconnect_0_sdram_0_s1_chipselect),                               //                                         .chipselect
		.seven_seg_pio_avalon_slave_0_address                (mm_interconnect_0_seven_seg_pio_avalon_slave_0_address),                //             seven_seg_pio_avalon_slave_0.address
		.seven_seg_pio_avalon_slave_0_write                  (mm_interconnect_0_seven_seg_pio_avalon_slave_0_write),                  //                                         .write
		.seven_seg_pio_avalon_slave_0_read                   (mm_interconnect_0_seven_seg_pio_avalon_slave_0_read),                   //                                         .read
		.seven_seg_pio_avalon_slave_0_readdata               (mm_interconnect_0_seven_seg_pio_avalon_slave_0_readdata),               //                                         .readdata
		.seven_seg_pio_avalon_slave_0_writedata              (mm_interconnect_0_seven_seg_pio_avalon_slave_0_writedata),              //                                         .writedata
		.seven_seg_pio_avalon_slave_0_chipselect             (mm_interconnect_0_seven_seg_pio_avalon_slave_0_chipselect),             //                                         .chipselect
		.spi_master_s1_address                               (mm_interconnect_0_spi_master_s1_address),                               //                            spi_master_s1.address
		.spi_master_s1_write                                 (mm_interconnect_0_spi_master_s1_write),                                 //                                         .write
		.spi_master_s1_read                                  (mm_interconnect_0_spi_master_s1_read),                                  //                                         .read
		.spi_master_s1_readdata                              (mm_interconnect_0_spi_master_s1_readdata),                              //                                         .readdata
		.spi_master_s1_writedata                             (mm_interconnect_0_spi_master_s1_writedata),                             //                                         .writedata
		.spi_master_s1_chipselect                            (mm_interconnect_0_spi_master_s1_chipselect),                            //                                         .chipselect
		.stimulus_in_s1_address                              (mm_interconnect_0_stimulus_in_s1_address),                              //                           stimulus_in_s1.address
		.stimulus_in_s1_write                                (mm_interconnect_0_stimulus_in_s1_write),                                //                                         .write
		.stimulus_in_s1_readdata                             (mm_interconnect_0_stimulus_in_s1_readdata),                             //                                         .readdata
		.stimulus_in_s1_writedata                            (mm_interconnect_0_stimulus_in_s1_writedata),                            //                                         .writedata
		.stimulus_in_s1_chipselect                           (mm_interconnect_0_stimulus_in_s1_chipselect),                           //                                         .chipselect
		.switch_pio_s1_address                               (mm_interconnect_0_switch_pio_s1_address),                               //                            switch_pio_s1.address
		.switch_pio_s1_readdata                              (mm_interconnect_0_switch_pio_s1_readdata),                              //                                         .readdata
		.sysid_qsys_0_control_slave_address                  (mm_interconnect_0_sysid_qsys_0_control_slave_address),                  //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                 (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),                 //                                         .readdata
		.system_timer_s1_address                             (mm_interconnect_0_system_timer_s1_address),                             //                          system_timer_s1.address
		.system_timer_s1_write                               (mm_interconnect_0_system_timer_s1_write),                               //                                         .write
		.system_timer_s1_readdata                            (mm_interconnect_0_system_timer_s1_readdata),                            //                                         .readdata
		.system_timer_s1_writedata                           (mm_interconnect_0_system_timer_s1_writedata),                           //                                         .writedata
		.system_timer_s1_chipselect                          (mm_interconnect_0_system_timer_s1_chipselect),                          //                                         .chipselect
		.timer_0_s1_address                                  (mm_interconnect_0_timer_0_s1_address),                                  //                               timer_0_s1.address
		.timer_0_s1_write                                    (mm_interconnect_0_timer_0_s1_write),                                    //                                         .write
		.timer_0_s1_readdata                                 (mm_interconnect_0_timer_0_s1_readdata),                                 //                                         .readdata
		.timer_0_s1_writedata                                (mm_interconnect_0_timer_0_s1_writedata),                                //                                         .writedata
		.timer_0_s1_chipselect                               (mm_interconnect_0_timer_0_s1_chipselect),                               //                                         .chipselect
		.uart_s1_address                                     (mm_interconnect_0_uart_s1_address),                                     //                                  uart_s1.address
		.uart_s1_write                                       (mm_interconnect_0_uart_s1_write),                                       //                                         .write
		.uart_s1_read                                        (mm_interconnect_0_uart_s1_read),                                        //                                         .read
		.uart_s1_readdata                                    (mm_interconnect_0_uart_s1_readdata),                                    //                                         .readdata
		.uart_s1_writedata                                   (mm_interconnect_0_uart_s1_writedata),                                   //                                         .writedata
		.uart_s1_begintransfer                               (mm_interconnect_0_uart_s1_begintransfer),                               //                                         .begintransfer
		.uart_s1_chipselect                                  (mm_interconnect_0_uart_s1_chipselect)                                   //                                         .chipselect
	);

	QD1_irq_mapper irq_mapper (
		.clk           (altpll_0_c2_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_0_c2_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_50_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
